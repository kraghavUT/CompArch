enum logic[4:0] { 
    ADD = 0,
    ADDI = 1,
    SUB = 2,
    SUBI = 3,
    MUL = 4,
    DIV = 5,
    AND = 6,
    OR = 7,
    XOR = 8,
    NOT = 9,
    SHFTR = 10,
    SHFTRI = 11,
    SHFTL = 12,
    SHFTLI = 13,
    BR = 14,
    BRR_R = 15,
    BRR_L = 16, 
    BRNZ = 17,
    CALL = 18,
    RETURN = 19,
    BRGT = 20,
    HALT = 31,
    MOV_MR = 21,
    MOV_RR = 22,
    MOV_RL = 23,
    MOV_RM = 24,
    ADDF = 25,
    SUBF = 26,
    MULF = 27,
    DIVF = 28,
    IN = 29,
    OUT = 30
} opcode_e;
